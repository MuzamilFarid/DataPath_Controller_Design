module control_fsm (
 
 input clk,
 input rst,
 





);






endmodule