module top_gcd ();

input wire clk,
input wire rst,




endmodule